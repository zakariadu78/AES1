library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library lib_aes;
library lib_rtl;
use lib_AES.state_definition_package.all;



entity Sbox_Inv_tb is 
end entity Sbox_Inv_tb; 


architecture Sbox_Inv_tb_arch of Sbox_Inv_tb is 
    component Sbox_Inv
    port (
    data_i  : in bit8; 
    data_o  : out bit8
    );
    end component;

signal data_i_s : bit8; 
signal data_o_s : bit8; 

begin 
    DUT : Sbox_Inv
        port map 
        (
            data_i => data_i_s,
            data_o => data_o_s
        );

P0 : process 
    begin 
        data_i_s <= x"00";
        wait for 10 ns; 
        data_i_s <= x"01";
        wait for 10 ns; 
        data_i_s <= x"02";
        wait for 10 ns; 
        data_i_s <= x"03";
        wait for 10 ns; 
        data_i_s <= x"04";
        wait for 10 ns; 
        data_i_s <= x"05";
        wait for 10 ns; 
        data_i_s <= x"06";
        wait for 10 ns; 
        data_i_s <= x"07";
        wait for 10 ns; 
        data_i_s <= x"08";
        wait for 10 ns; 
        data_i_s <= x"09";
        wait for 10 ns; 
        data_i_s <= x"10";
        wait for 10 ns; 
        data_i_s <= x"0A";
        wait for 10 ns; 
        data_i_s <= x"0B";
        wait for 10 ns;
        data_i_s <= x"0C";
        wait for 10 ns;  
        data_i_s <= x"0D";
        wait for 10 ns; 
        data_i_s <= x"0E";
        wait for 10 ns; 

        data_i_s <= x"10";
        wait for 10 ns; 
        data_i_s <= x"11";
        wait for 10 ns; 
        data_i_s <= x"12";
        wait for 10 ns; 
        data_i_s <= x"13";
        wait for 10 ns; 
        data_i_s <= x"14";
        wait for 10 ns; 
        data_i_s <= x"15";
        wait for 10 ns; 
        data_i_s <= x"16";
        wait for 10 ns; 
        data_i_s <= x"17";
        wait for 10 ns; 
        data_i_s <= x"18";
        wait for 10 ns; 
        data_i_s <= x"19";
        wait for 10 ns; 
        data_i_s <= x"1A";
        wait for 10 ns; 
        data_i_s <= x"1B";
        wait for 10 ns;
        data_i_s <= x"1C";
        wait for 10 ns;  
        data_i_s <= x"1D";
        wait for 10 ns; 
        data_i_s <= x"1E";
        wait for 10 ns; 
        
        data_i_s <= x"20";
        wait for 10 ns; 
        data_i_s <= x"21";
        wait for 10 ns; 
        data_i_s <= x"22";
        wait for 10 ns; 
        data_i_s <= x"23";
        wait for 10 ns; 
        data_i_s <= x"24";
        wait for 10 ns; 
        data_i_s <= x"25";
        wait for 10 ns; 
        data_i_s <= x"26";
        wait for 10 ns; 
        data_i_s <= x"27";
        wait for 10 ns; 
        data_i_s <= x"28";
        wait for 10 ns; 
        data_i_s <= x"29";
        wait for 10 ns; 
        data_i_s <= x"2A";
        wait for 10 ns; 
        data_i_s <= x"2B";
        wait for 10 ns;
        data_i_s <= x"2C";
        wait for 10 ns;  
        data_i_s <= x"2D";
        wait for 10 ns; 
        data_i_s <= x"2E";
        wait for 10 ns;

        data_i_s <= x"30";
        wait for 10 ns; 
        data_i_s <= x"31";
        wait for 10 ns; 
        data_i_s <= x"32";
        wait for 10 ns; 
        data_i_s <= x"33";
        wait for 10 ns; 
        data_i_s <= x"34";
        wait for 10 ns; 
        data_i_s <= x"35";
        wait for 10 ns; 
        data_i_s <= x"36";
        wait for 10 ns; 
        data_i_s <= x"37";
        wait for 10 ns; 
        data_i_s <= x"38";
        wait for 10 ns; 
        data_i_s <= x"39";
        wait for 10 ns; 
        data_i_s <= x"3A";
        wait for 10 ns; 
        data_i_s <= x"3B";
        wait for 10 ns;
        data_i_s <= x"3C";
        wait for 10 ns;  
        data_i_s <= x"3D";
        wait for 10 ns; 
        data_i_s <= x"3E";
        wait for 10 ns;

        data_i_s <= x"40";
        wait for 10 ns; 
        data_i_s <= x"41";
        wait for 10 ns; 
        data_i_s <= x"42";
        wait for 10 ns; 
        data_i_s <= x"43";
        wait for 10 ns; 
        data_i_s <= x"44";
        wait for 10 ns; 
        data_i_s <= x"45";
        wait for 10 ns; 
        data_i_s <= x"46";
        wait for 10 ns; 
        data_i_s <= x"47";
        wait for 10 ns; 
        data_i_s <= x"48";
        wait for 10 ns; 
        data_i_s <= x"49";
        wait for 10 ns; 
        data_i_s <= x"4A";
        wait for 10 ns; 
        data_i_s <= x"4B";
        wait for 10 ns;
        data_i_s <= x"4C";
        wait for 10 ns;  
        data_i_s <= x"4D";
        wait for 10 ns; 
        data_i_s <= x"4E";
        wait for 10 ns;
         
        data_i_s <= x"50";
        wait for 10 ns; 
        data_i_s <= x"51";
        wait for 10 ns; 
        data_i_s <= x"52";
        wait for 10 ns; 
        data_i_s <= x"53";
        wait for 10 ns; 
        data_i_s <= x"54";
        wait for 10 ns; 
        data_i_s <= x"55";
        wait for 10 ns; 
        data_i_s <= x"56";
        wait for 10 ns; 
        data_i_s <= x"57";
        wait for 10 ns; 
        data_i_s <= x"58";
        wait for 10 ns; 
        data_i_s <= x"59";
        wait for 10 ns; 
        data_i_s <= x"5A";
        wait for 10 ns; 
        data_i_s <= x"5B";
        wait for 10 ns;
        data_i_s <= x"5C";
        wait for 10 ns;  
        data_i_s <= x"5D";
        wait for 10 ns; 
        data_i_s <= x"5E";
        wait for 10 ns;

        data_i_s <= x"60";
        wait for 10 ns; 
        data_i_s <= x"61";
        wait for 10 ns; 
        data_i_s <= x"62";
        wait for 10 ns; 
        data_i_s <= x"63";
        wait for 10 ns; 
        data_i_s <= x"64";
        wait for 10 ns; 
        data_i_s <= x"65";
        wait for 10 ns; 
        data_i_s <= x"66";
        wait for 10 ns; 
        data_i_s <= x"67";
        wait for 10 ns; 
        data_i_s <= x"68";
        wait for 10 ns; 
        data_i_s <= x"69";
        wait for 10 ns; 
        data_i_s <= x"6A";
        wait for 10 ns; 
        data_i_s <= x"6B";
        wait for 10 ns;
        data_i_s <= x"6C";
        wait for 10 ns;  
        data_i_s <= x"6D";
        wait for 10 ns; 
        data_i_s <= x"6E";
        wait for 10 ns;

        data_i_s <= x"70";
        wait for 10 ns; 
        data_i_s <= x"71";
        wait for 10 ns; 
        data_i_s <= x"72";
        wait for 10 ns; 
        data_i_s <= x"73";
        wait for 10 ns; 
        data_i_s <= x"74";
        wait for 10 ns; 
        data_i_s <= x"75";
        wait for 10 ns; 
        data_i_s <= x"76";
        wait for 10 ns; 
        data_i_s <= x"77";
        wait for 10 ns; 
        data_i_s <= x"78";
        wait for 10 ns; 
        data_i_s <= x"79";
        wait for 10 ns; 
        data_i_s <= x"7A";
        wait for 10 ns; 
        data_i_s <= x"7B";
        wait for 10 ns;
        data_i_s <= x"7C";
        wait for 10 ns;  
        data_i_s <= x"7D";
        wait for 10 ns; 
        data_i_s <= x"7E";
        wait for 10 ns;

        data_i_s <= x"80";
        wait for 10 ns; 
        data_i_s <= x"81";
        wait for 10 ns; 
        data_i_s <= x"82";
        wait for 10 ns; 
        data_i_s <= x"83";
        wait for 10 ns; 
        data_i_s <= x"84";
        wait for 10 ns; 
        data_i_s <= x"85";
        wait for 10 ns; 
        data_i_s <= x"86";
        wait for 10 ns; 
        data_i_s <= x"87";
        wait for 10 ns; 
        data_i_s <= x"88";
        wait for 10 ns; 
        data_i_s <= x"89";
        wait for 10 ns; 
        data_i_s <= x"8A";
        wait for 10 ns; 
        data_i_s <= x"8B";
        wait for 10 ns;
        data_i_s <= x"8C";
        wait for 10 ns;  
        data_i_s <= x"8D";
        wait for 10 ns; 
        data_i_s <= x"8E";
        wait for 10 ns;

        data_i_s <= x"90";
        wait for 10 ns; 
        data_i_s <= x"91";
        wait for 10 ns; 
        data_i_s <= x"92";
        wait for 10 ns; 
        data_i_s <= x"93";
        wait for 10 ns; 
        data_i_s <= x"94";
        wait for 10 ns; 
        data_i_s <= x"95";
        wait for 10 ns; 
        data_i_s <= x"96";
        wait for 10 ns; 
        data_i_s <= x"97";
        wait for 10 ns; 
        data_i_s <= x"98";
        wait for 10 ns; 
        data_i_s <= x"99";
        wait for 10 ns; 
        data_i_s <= x"9A";
        wait for 10 ns; 
        data_i_s <= x"9B";
        wait for 10 ns;
        data_i_s <= x"9C";
        wait for 10 ns;  
        data_i_s <= x"9D";
        wait for 10 ns; 
        data_i_s <= x"9E";
        wait for 10 ns;

end process P0;
end architecture;