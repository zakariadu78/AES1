-- Pas nécessaire, testé directement sur l'AES Global