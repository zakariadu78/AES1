LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
LIBRARY lib_rtl;
LIBRARY lib_aes;
USE lib_aes.state_definition_package.ALL;

ENTITY Sbox_Inv_tb IS
END ENTITY Sbox_Inv_tb;
ARCHITECTURE Sbox_Inv_tb_arch OF Sbox_Inv_tb IS
    COMPONENT Sbox_Inv
        PORT (
            data_i : IN bit8;
            data_o : OUT bit8
        );
    END COMPONENT;

    SIGNAL data_i_s : bit8;
    SIGNAL data_o_s : bit8;

BEGIN
    DUT : Sbox_Inv
    PORT MAP
    (
        data_i => data_i_s,
        data_o => data_o_s
    );

    P0 : PROCESS
    BEGIN
        data_i_s <= x"00";
        WAIT FOR 10 ns;
        data_i_s <= x"01";
        WAIT FOR 10 ns;
        data_i_s <= x"02";
        WAIT FOR 10 ns;
        data_i_s <= x"03";
        WAIT FOR 10 ns;
        data_i_s <= x"04";
        WAIT FOR 10 ns;
        data_i_s <= x"05";
        WAIT FOR 10 ns;
        data_i_s <= x"06";
        WAIT FOR 10 ns;
        data_i_s <= x"07";
        WAIT FOR 10 ns;
        data_i_s <= x"08";
        WAIT FOR 10 ns;
        data_i_s <= x"09";
        WAIT FOR 10 ns;
        data_i_s <= x"10";
        WAIT FOR 10 ns;
        data_i_s <= x"0A";
        WAIT FOR 10 ns;
        data_i_s <= x"0B";
        WAIT FOR 10 ns;
        data_i_s <= x"0C";
        WAIT FOR 10 ns;
        data_i_s <= x"0D";
        WAIT FOR 10 ns;
        data_i_s <= x"0E";
        WAIT FOR 10 ns;

        data_i_s <= x"10";
        WAIT FOR 10 ns;
        data_i_s <= x"11";
        WAIT FOR 10 ns;
        data_i_s <= x"12";
        WAIT FOR 10 ns;
        data_i_s <= x"13";
        WAIT FOR 10 ns;
        data_i_s <= x"14";
        WAIT FOR 10 ns;
        data_i_s <= x"15";
        WAIT FOR 10 ns;
        data_i_s <= x"16";
        WAIT FOR 10 ns;
        data_i_s <= x"17";
        WAIT FOR 10 ns;
        data_i_s <= x"18";
        WAIT FOR 10 ns;
        data_i_s <= x"19";
        WAIT FOR 10 ns;
        data_i_s <= x"1A";
        WAIT FOR 10 ns;
        data_i_s <= x"1B";
        WAIT FOR 10 ns;
        data_i_s <= x"1C";
        WAIT FOR 10 ns;
        data_i_s <= x"1D";
        WAIT FOR 10 ns;
        data_i_s <= x"1E";
        WAIT FOR 10 ns;

        data_i_s <= x"20";
        WAIT FOR 10 ns;
        data_i_s <= x"21";
        WAIT FOR 10 ns;
        data_i_s <= x"22";
        WAIT FOR 10 ns;
        data_i_s <= x"23";
        WAIT FOR 10 ns;
        data_i_s <= x"24";
        WAIT FOR 10 ns;
        data_i_s <= x"25";
        WAIT FOR 10 ns;
        data_i_s <= x"26";
        WAIT FOR 10 ns;
        data_i_s <= x"27";
        WAIT FOR 10 ns;
        data_i_s <= x"28";
        WAIT FOR 10 ns;
        data_i_s <= x"29";
        WAIT FOR 10 ns;
        data_i_s <= x"2A";
        WAIT FOR 10 ns;
        data_i_s <= x"2B";
        WAIT FOR 10 ns;
        data_i_s <= x"2C";
        WAIT FOR 10 ns;
        data_i_s <= x"2D";
        WAIT FOR 10 ns;
        data_i_s <= x"2E";
        WAIT FOR 10 ns;

        data_i_s <= x"30";
        WAIT FOR 10 ns;
        data_i_s <= x"31";
        WAIT FOR 10 ns;
        data_i_s <= x"32";
        WAIT FOR 10 ns;
        data_i_s <= x"33";
        WAIT FOR 10 ns;
        data_i_s <= x"34";
        WAIT FOR 10 ns;
        data_i_s <= x"35";
        WAIT FOR 10 ns;
        data_i_s <= x"36";
        WAIT FOR 10 ns;
        data_i_s <= x"37";
        WAIT FOR 10 ns;
        data_i_s <= x"38";
        WAIT FOR 10 ns;
        data_i_s <= x"39";
        WAIT FOR 10 ns;
        data_i_s <= x"3A";
        WAIT FOR 10 ns;
        data_i_s <= x"3B";
        WAIT FOR 10 ns;
        data_i_s <= x"3C";
        WAIT FOR 10 ns;
        data_i_s <= x"3D";
        WAIT FOR 10 ns;
        data_i_s <= x"3E";
        WAIT FOR 10 ns;

        data_i_s <= x"40";
        WAIT FOR 10 ns;
        data_i_s <= x"41";
        WAIT FOR 10 ns;
        data_i_s <= x"42";
        WAIT FOR 10 ns;
        data_i_s <= x"43";
        WAIT FOR 10 ns;
        data_i_s <= x"44";
        WAIT FOR 10 ns;
        data_i_s <= x"45";
        WAIT FOR 10 ns;
        data_i_s <= x"46";
        WAIT FOR 10 ns;
        data_i_s <= x"47";
        WAIT FOR 10 ns;
        data_i_s <= x"48";
        WAIT FOR 10 ns;
        data_i_s <= x"49";
        WAIT FOR 10 ns;
        data_i_s <= x"4A";
        WAIT FOR 10 ns;
        data_i_s <= x"4B";
        WAIT FOR 10 ns;
        data_i_s <= x"4C";
        WAIT FOR 10 ns;
        data_i_s <= x"4D";
        WAIT FOR 10 ns;
        data_i_s <= x"4E";
        WAIT FOR 10 ns;

        data_i_s <= x"50";
        WAIT FOR 10 ns;
        data_i_s <= x"51";
        WAIT FOR 10 ns;
        data_i_s <= x"52";
        WAIT FOR 10 ns;
        data_i_s <= x"53";
        WAIT FOR 10 ns;
        data_i_s <= x"54";
        WAIT FOR 10 ns;
        data_i_s <= x"55";
        WAIT FOR 10 ns;
        data_i_s <= x"56";
        WAIT FOR 10 ns;
        data_i_s <= x"57";
        WAIT FOR 10 ns;
        data_i_s <= x"58";
        WAIT FOR 10 ns;
        data_i_s <= x"59";
        WAIT FOR 10 ns;
        data_i_s <= x"5A";
        WAIT FOR 10 ns;
        data_i_s <= x"5B";
        WAIT FOR 10 ns;
        data_i_s <= x"5C";
        WAIT FOR 10 ns;
        data_i_s <= x"5D";
        WAIT FOR 10 ns;
        data_i_s <= x"5E";
        WAIT FOR 10 ns;

        data_i_s <= x"60";
        WAIT FOR 10 ns;
        data_i_s <= x"61";
        WAIT FOR 10 ns;
        data_i_s <= x"62";
        WAIT FOR 10 ns;
        data_i_s <= x"63";
        WAIT FOR 10 ns;
        data_i_s <= x"64";
        WAIT FOR 10 ns;
        data_i_s <= x"65";
        WAIT FOR 10 ns;
        data_i_s <= x"66";
        WAIT FOR 10 ns;
        data_i_s <= x"67";
        WAIT FOR 10 ns;
        data_i_s <= x"68";
        WAIT FOR 10 ns;
        data_i_s <= x"69";
        WAIT FOR 10 ns;
        data_i_s <= x"6A";
        WAIT FOR 10 ns;
        data_i_s <= x"6B";
        WAIT FOR 10 ns;
        data_i_s <= x"6C";
        WAIT FOR 10 ns;
        data_i_s <= x"6D";
        WAIT FOR 10 ns;
        data_i_s <= x"6E";
        WAIT FOR 10 ns;

        data_i_s <= x"70";
        WAIT FOR 10 ns;
        data_i_s <= x"71";
        WAIT FOR 10 ns;
        data_i_s <= x"72";
        WAIT FOR 10 ns;
        data_i_s <= x"73";
        WAIT FOR 10 ns;
        data_i_s <= x"74";
        WAIT FOR 10 ns;
        data_i_s <= x"75";
        WAIT FOR 10 ns;
        data_i_s <= x"76";
        WAIT FOR 10 ns;
        data_i_s <= x"77";
        WAIT FOR 10 ns;
        data_i_s <= x"78";
        WAIT FOR 10 ns;
        data_i_s <= x"79";
        WAIT FOR 10 ns;
        data_i_s <= x"7A";
        WAIT FOR 10 ns;
        data_i_s <= x"7B";
        WAIT FOR 10 ns;
        data_i_s <= x"7C";
        WAIT FOR 10 ns;
        data_i_s <= x"7D";
        WAIT FOR 10 ns;
        data_i_s <= x"7E";
        WAIT FOR 10 ns;

        data_i_s <= x"80";
        WAIT FOR 10 ns;
        data_i_s <= x"81";
        WAIT FOR 10 ns;
        data_i_s <= x"82";
        WAIT FOR 10 ns;
        data_i_s <= x"83";
        WAIT FOR 10 ns;
        data_i_s <= x"84";
        WAIT FOR 10 ns;
        data_i_s <= x"85";
        WAIT FOR 10 ns;
        data_i_s <= x"86";
        WAIT FOR 10 ns;
        data_i_s <= x"87";
        WAIT FOR 10 ns;
        data_i_s <= x"88";
        WAIT FOR 10 ns;
        data_i_s <= x"89";
        WAIT FOR 10 ns;
        data_i_s <= x"8A";
        WAIT FOR 10 ns;
        data_i_s <= x"8B";
        WAIT FOR 10 ns;
        data_i_s <= x"8C";
        WAIT FOR 10 ns;
        data_i_s <= x"8D";
        WAIT FOR 10 ns;
        data_i_s <= x"8E";
        WAIT FOR 10 ns;

        data_i_s <= x"90";
        WAIT FOR 10 ns;
        data_i_s <= x"91";
        WAIT FOR 10 ns;
        data_i_s <= x"92";
        WAIT FOR 10 ns;
        data_i_s <= x"93";
        WAIT FOR 10 ns;
        data_i_s <= x"94";
        WAIT FOR 10 ns;
        data_i_s <= x"95";
        WAIT FOR 10 ns;
        data_i_s <= x"96";
        WAIT FOR 10 ns;
        data_i_s <= x"97";
        WAIT FOR 10 ns;
        data_i_s <= x"98";
        WAIT FOR 10 ns;
        data_i_s <= x"99";
        WAIT FOR 10 ns;
        data_i_s <= x"9A";
        WAIT FOR 10 ns;
        data_i_s <= x"9B";
        WAIT FOR 10 ns;
        data_i_s <= x"9C";
        WAIT FOR 10 ns;
        data_i_s <= x"9D";
        WAIT FOR 10 ns;
        data_i_s <= x"9E";
        WAIT FOR 10 ns;

    END PROCESS P0;
END ARCHITECTURE;