library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library lib_rtl;
use lib_rtl.state_definition_package.all;



entity Sbox_tb is 
end entity Sbox_tb; 


architecture Sbox_tb_arch of Sbox_tb is 
    component Sbox_tb
    port (
    data_i  : in bit8; 
    data_o  : out bit8
    );
    end component;

signal data_i_s : bit8; 
signal data_o_s : bit8; 

begin 
    DUT : Sbox
        port map 
        (
            data_i => data_i_s,
            data_o => data_o_s
        );

P0 : process 
    begin 
        data_i <= x"00";
        wait for 10ns; 
        data_i <= x"01";
        wait for 10ns; 
        data_i <= x"02";
        wait for 10ns; 
        data_i <= x"03";
        wait for 10ns; 
        data_i <= x"04";
        wait for 10ns; 
        data_i <= x"05";
        wait for 10ns; 
        data_i <= x"06";
        wait for 10ns; 
        data_i <= x"07";
        wait for 10ns; 
        data_i <= x"08";
        wait for 10ns; 
        data_i <= x"09";
        wait for 10ns; 
        data_i <= x"10";
        wait for 10ns; 
        data_i <= x"0A";
        wait for 10ns; 
        data_i <= x"0B";
        wait for 10ns;
        data_i <= x"0C";
        wait for 10ns;  
        data_i <= x"0D";
        wait for 10ns; 
        data_i <= x"0E";
        wait for 10ns; 

        data_i <= x"10";
        wait for 10ns; 
        data_i <= x"11";
        wait for 10ns; 
        data_i <= x"12";
        wait for 10ns; 
        data_i <= x"13";
        wait for 10ns; 
        data_i <= x"14";
        wait for 10ns; 
        data_i <= x"15";
        wait for 10ns; 
        data_i <= x"16";
        wait for 10ns; 
        data_i <= x"17";
        wait for 10ns; 
        data_i <= x"18";
        wait for 10ns; 
        data_i <= x"19";
        wait for 10ns; 
        data_i <= x"1A";
        wait for 10ns; 
        data_i <= x"1B";
        wait for 10ns;
        data_i <= x"1C";
        wait for 10ns;  
        data_i <= x"1D";
        wait for 10ns; 
        data_i <= x"1E";
        wait for 10ns; 
        
        data_i <= x"20";
        wait for 10ns; 
        data_i <= x"21";
        wait for 10ns; 
        data_i <= x"22";
        wait for 10ns; 
        data_i <= x"23";
        wait for 10ns; 
        data_i <= x"24";
        wait for 10ns; 
        data_i <= x"25";
        wait for 10ns; 
        data_i <= x"26";
        wait for 10ns; 
        data_i <= x"27";
        wait for 10ns; 
        data_i <= x"28";
        wait for 10ns; 
        data_i <= x"29";
        wait for 10ns; 
        data_i <= x"2A";
        wait for 10ns; 
        data_i <= x"2B";
        wait for 10ns;
        data_i <= x"2C";
        wait for 10ns;  
        data_i <= x"2D";
        wait for 10ns; 
        data_i <= x"2E";
        wait for 10ns;

        data_i <= x"30";
        wait for 10ns; 
        data_i <= x"31";
        wait for 10ns; 
        data_i <= x"32";
        wait for 10ns; 
        data_i <= x"33";
        wait for 10ns; 
        data_i <= x"34";
        wait for 10ns; 
        data_i <= x"35";
        wait for 10ns; 
        data_i <= x"36";
        wait for 10ns; 
        data_i <= x"37";
        wait for 10ns; 
        data_i <= x"38";
        wait for 10ns; 
        data_i <= x"39";
        wait for 10ns; 
        data_i <= x"3A";
        wait for 10ns; 
        data_i <= x"3B";
        wait for 10ns;
        data_i <= x"3C";
        wait for 10ns;  
        data_i <= x"3D";
        wait for 10ns; 
        data_i <= x"3E";
        wait for 10ns;

        data_i <= x"40";
        wait for 10ns; 
        data_i <= x"41";
        wait for 10ns; 
        data_i <= x"42";
        wait for 10ns; 
        data_i <= x"43";
        wait for 10ns; 
        data_i <= x"44";
        wait for 10ns; 
        data_i <= x"45";
        wait for 10ns; 
        data_i <= x"46";
        wait for 10ns; 
        data_i <= x"47";
        wait for 10ns; 
        data_i <= x"48";
        wait for 10ns; 
        data_i <= x"49";
        wait for 10ns; 
        data_i <= x"4A";
        wait for 10ns; 
        data_i <= x"4B";
        wait for 10ns;
        data_i <= x"4C";
        wait for 10ns;  
        data_i <= x"4D";
        wait for 10ns; 
        data_i <= x"4E";
        wait for 10ns;
         
        data_i <= x"50";
        wait for 10ns; 
        data_i <= x"51";
        wait for 10ns; 
        data_i <= x"52";
        wait for 10ns; 
        data_i <= x"53";
        wait for 10ns; 
        data_i <= x"54";
        wait for 10ns; 
        data_i <= x"55";
        wait for 10ns; 
        data_i <= x"56";
        wait for 10ns; 
        data_i <= x"57";
        wait for 10ns; 
        data_i <= x"58";
        wait for 10ns; 
        data_i <= x"59";
        wait for 10ns; 
        data_i <= x"5A";
        wait for 10ns; 
        data_i <= x"5B";
        wait for 10ns;
        data_i <= x"5C";
        wait for 10ns;  
        data_i <= x"5D";
        wait for 10ns; 
        data_i <= x"5E";
        wait for 10ns;

        data_i <= x"60";
        wait for 10ns; 
        data_i <= x"61";
        wait for 10ns; 
        data_i <= x"62";
        wait for 10ns; 
        data_i <= x"63";
        wait for 10ns; 
        data_i <= x"64";
        wait for 10ns; 
        data_i <= x"65";
        wait for 10ns; 
        data_i <= x"66";
        wait for 10ns; 
        data_i <= x"67";
        wait for 10ns; 
        data_i <= x"68";
        wait for 10ns; 
        data_i <= x"69";
        wait for 10ns; 
        data_i <= x"6A";
        wait for 10ns; 
        data_i <= x"6B";
        wait for 10ns;
        data_i <= x"6C";
        wait for 10ns;  
        data_i <= x"6D";
        wait for 10ns; 
        data_i <= x"6E";
        wait for 10ns;

        data_i <= x"70";
        wait for 10ns; 
        data_i <= x"71";
        wait for 10ns; 
        data_i <= x"72";
        wait for 10ns; 
        data_i <= x"73";
        wait for 10ns; 
        data_i <= x"74";
        wait for 10ns; 
        data_i <= x"75";
        wait for 10ns; 
        data_i <= x"76";
        wait for 10ns; 
        data_i <= x"77";
        wait for 10ns; 
        data_i <= x"78";
        wait for 10ns; 
        data_i <= x"79";
        wait for 10ns; 
        data_i <= x"7A";
        wait for 10ns; 
        data_i <= x"7B";
        wait for 10ns;
        data_i <= x"7C";
        wait for 10ns;  
        data_i <= x"7D";
        wait for 10ns; 
        data_i <= x"7E";
        wait for 10ns;

        data_i <= x"80";
        wait for 10ns; 
        data_i <= x"81";
        wait for 10ns; 
        data_i <= x"82";
        wait for 10ns; 
        data_i <= x"83";
        wait for 10ns; 
        data_i <= x"84";
        wait for 10ns; 
        data_i <= x"85";
        wait for 10ns; 
        data_i <= x"86";
        wait for 10ns; 
        data_i <= x"87";
        wait for 10ns; 
        data_i <= x"88";
        wait for 10ns; 
        data_i <= x"89";
        wait for 10ns; 
        data_i <= x"8A";
        wait for 10ns; 
        data_i <= x"8B";
        wait for 10ns;
        data_i <= x"8C";
        wait for 10ns;  
        data_i <= x"8D";
        wait for 10ns; 
        data_i <= x"8E";
        wait for 10ns;

        data_i <= x"90";
        wait for 10ns; 
        data_i <= x"91";
        wait for 10ns; 
        data_i <= x"92";
        wait for 10ns; 
        data_i <= x"93";
        wait for 10ns; 
        data_i <= x"94";
        wait for 10ns; 
        data_i <= x"95";
        wait for 10ns; 
        data_i <= x"96";
        wait for 10ns; 
        data_i <= x"97";
        wait for 10ns; 
        data_i <= x"98";
        wait for 10ns; 
        data_i <= x"99";
        wait for 10ns; 
        data_i <= x"9A";
        wait for 10ns; 
        data_i <= x"9B";
        wait for 10ns;
        data_i <= x"9C";
        wait for 10ns;  
        data_i <= x"9D";
        wait for 10ns; 
        data_i <= x"9E";
        wait for 10ns;

end process P0;
end architecture Sbox_tb_arch;